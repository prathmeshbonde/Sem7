
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity usr44 is
    Port ( Rst : in  STD_LOGIC;
           Clk : in  STD_LOGIC;
           Sin : in  STD_LOGIC;
           Pin : in  STD_LOGIC_VECTOR (3 downto 0);
           Mode : in  STD_LOGIC_VECTOR (1 downto 0);
           Sout : out  STD_LOGIC;
           Pout : out  STD_LOGIC_VECTOR (3 downto 0));
end usr44;

architecture usr44_arch of usr44 is

begin


end usr44_arch;

